library verilog;
use verilog.vl_types.all;
entity TestBenchRepair is
end TestBenchRepair;
