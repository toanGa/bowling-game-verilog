library verilog;
use verilog.vl_types.all;
entity TestLed is
end TestLed;
